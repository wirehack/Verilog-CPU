`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:48:46 10/19/2015 
// Design Name: 
// Module Name:    decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder(
    input x0,
    input x1,
    input x2,
    input x3,
    output a,
    output b,
    output c,
    output d,
    output e,
    output f,
    output g
    );
    reg a,b,c,d,e,f,g;
    always@*
    begin
        assign a=(!x3 && !x2 && !x1 && !x0) || (!x3 && !x2 && x1 && !x0) || (!x3 && !x2 && x1 && x0) || (!x3 && x2 && !x1 && x0) || (!x3 && x2 && x1 && !x0) || (!x3 && x2 && x1 && x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && !x0) || (x3 && x2 && !x1 && !x0) || (x3 && x2 && x1 && !x0) || (x3 && x2 && x1 && x0);
        assign b=(!x3 && !x2 && !x1 && !x0) || (!x3 && x2 && !x1 && !x0) || (!x3 && x2 && !x1 && x0) || (!x3 && x2 && x1 && !x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && !x0) || (x3 && !x2 && x1 && x0) || (x3 && x2 && !x1 && !x0) || (x3 && x2 && x1 && !x0) || (x3 && x2 && x1 && x0);
        assign c=(!x3 && !x2 && !x1 && !x0) || (!x3 && !x2 && x1 && !x0) || (!x3 && x2 && x1 && !x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && x1 && !x0) || (x3 && !x2 && x1 && x0) || (x3 && x2 && !x1 && !x0) || (x3 && x2 && !x1 && x0) || (x3 && x2 && x1 && !x0) || (x3 && x2 && x1 && x0);
        assign d=(!x3 && !x2 && !x1 && !x0) || (!x3 && !x2 && x1 && !x0) || (!x3 && !x2 && x1 && x0) || (!x3 && x2 && !x1 && x0) || (!x3 && x2 && x1 && !x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && x0) || (x3 && x2 && !x1 && !x0) || (x3 && x2 && !x1 && x0) || (x3 && x2 && x1 && !x0);
        assign e=(!x3 && !x2 && !x1 && !x0) || (!x3 && !x2 && !x1 && x0) || (!x3 && !x2 && x1 && x0) || (!x3 && x2 && !x1 && !x0) || (!x3 && x2 && !x1 && x0) || (!x3 && x2 && x1 && !x0) || (!x3 && x2 && x1 && x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && !x0) || (x3 && !x2 && x1 && x0) || (x3 && x2 && !x1 && x0);
        assign f=(!x3 && !x2 && !x1 && !x0) || (!x3 && !x2 && !x1 && x0) || (!x3 && !x2 && x1 && !x0) || (!x3 && !x2 && x1 && x0) || (!x3 && x2 && !x1 && !x0) || (!x3 && x2 && x1 && x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && !x0) || (x3 && x2 && !x1 && x0);
        assign g=(!x3 && !x2 && x1 && !x0) || (!x3 && !x2 && x1 && x0) || (!x3 && x2 && !x1 && !x0) || (!x3 && x2 && !x1 && x0) || (!x3 && x2 && x1 && !x0) || (x3 && !x2 && !x1 && !x0) || (x3 && !x2 && !x1 && x0) || (x3 && !x2 && x1 && !x0) || (x3 && !x2 && x1 && x0) || (x3 && x2 && !x1 && x0) || (x3 && x2 && x1 && !x0) || (x3 && x2 && x1 && x0);
    end
endmodule
